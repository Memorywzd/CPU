//指令寄存器，存储要执行的指令
//注意：该寄存器是时钟的下降沿有效

module ir(din,clk,rst,irload,dout);

endmodule