//R通用寄存器，用来存放第二个操作数

module r(din, clk, rst,rload, dout);

endmodule
