//AC通用寄存器，存储第一个操作数

module ac(din, clk, rst,acload, dout);

endmodule
