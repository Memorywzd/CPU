//标志寄存器

module z(din,clk,rst, zload,dout);

endmodule