//算术逻辑单元

module alu(alus,ac, bus, dout);


endmodule
