//数据暂存器,处理双字节指令时使用，用来存储低八位的地址或数值

module tr(din, clk,rst, trload, dout);

endmodule