//将cpu组件实例化后定义cpu组件

module cpu_obj(data_in,clk_quick,clk_slow,clk_delay,rst,SW_choose,A1,cpustate,addr,data_out,acdbus,rdbus,...... ,clr);


endmodule
