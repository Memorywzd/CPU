//数据寄存器，存放双指令中低8位指向地址的存放值

module dr(din, clk,rst, drload, dout);

endmodule